module Fourth_les(
input wire [3:0] SW, // ????????????? ????? (??????? A)
output wire [4:0] LEDR // ?????????? ?????: sum[3:0], cout
);
wire [3:0] a = SW[3:0];
wire [3:0] b = 4'd7; // 
wire cin = 1'b0; // 
adder_4bit DUT(
.a(a),
.b(b),
.cin(cin),
.sum(LEDR[3:0]),
.cout(LEDR[4])
);
endmodule
