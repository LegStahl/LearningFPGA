module memory();



endmodule