

// Определение модуля и его портов ввода/вывода
module universal_shift_reg (
    // ----------- Входные порты -----------
    input wire         clk,           // Тактовый сигнал. Все синхронные операции выполняются по его положительному фронту.
    input wire         rst_n,         // Асинхронный сброс, активный уровень - низкий ('0'). При сбросе выход обнуляется.
    input wire   [1:0] select,        // Управляющий сигнал для выбора режима работы регистра.
    input wire   [3:0] p_din,         // 4-битная шина для параллельной загрузки данных.
    input wire         s_left_din,    // Входной бит для операции сдвига влево (загружается в LSB).
    input wire         s_right_din,   // Входной бит для операции сдвига вправо (загружается в MSB).

    // ----------- Выходные порты ----------
    output reg   [3:0] p_dout         // 4-битный выход регистра. Объявлен как 'reg', так как его значение
                                      // присваивается внутри процедурного блока 'always'.
);

    // Основной процедурный блок, описывающий поведение регистра.
    // Блок чувствителен к положительному фронту тактового сигнала (posedge clk)
    // и к отрицательному уровню сигнала сброса (negedge rst_n).
    // Это стандартный шаблон для описания синхронной логики с асинхронным сбросом.
    always @(posedge clk or negedge rst_n) begin
        // --- Логика асинхронного сброса ---
        // Если сигнал сброса 'rst_n' находится в активном (низком) состоянии,
        // выходное значение регистра немедленно обнуляется,
        // игнорируя тактовый сигнал и другие входы.
        if (!rst_n) begin
            p_dout <= 4'b0000; // Используется неблокирующее присваивание '<=' для регистровой логики.
        end
        // --- Синхронная логика работы ---
        // Если сброс неактивен, модуль работает в синхронном режиме.
        // Все изменения происходят только по положительному фронту 'clk'.
        else begin
            // Конструкция 'case' используется для выбора операции в зависимости
            // от значения управляющего сигнала 'select'.
            case (select)
                // Режим 2'b00: Хранение (Hold)
                // Выходное значение регистра не меняется, сохраняя свое предыдущее состояние.
                2'b00: begin
                    p_dout <= p_dout;
                end

                // Режим 2'b01: Логический сдвиг вправо (Shift Right)
                // Старший бит (MSB) p_dout[3] принимает значение с входа s_right_din.
                // Остальные биты [2:0] сдвигаются на одну позицию вправо.
                // Младший бит (LSB) p_dout[0] отбрасывается.
                // Пример: если p_dout = 1011 и s_right_din = 0, новым значением будет 0101.
                2'b01: begin
                    p_dout <= {s_right_din, p_dout[3:1]}; // Оператор конкатенации {} для формирования нового значения.
                end

                // Режим 2'b10: Логический сдвиг влево (Shift Left)
                // Младший бит (LSB) p_dout[0] принимает значение с входа s_left_din.
                // Остальные биты [3:1] сдвигаются на одну позицию влево.
                // Старший бит (MSB) p_dout[3] отбрасывается.
                // Пример: если p_dout = 1011 и s_left_din = 0, новым значением будет 0110.
                2'b10: begin
                    p_dout <= {p_dout[2:0], s_left_din};
                end

                // Режим 2'b11: Параллельная загрузка (Parallel Load)
                // Регистр полностью загружает 4-битное значение с входа p_din.
                2'b11: begin
                    p_dout <= p_din;
                end

                // Ветвь 'default': на случай неопределенных или 'x'/'z' состояний на 'select'.
                // Чтобы избежать неявного создания "защелок" (latches) при синтезе,
                // рекомендуется всегда определять поведение для всех возможных случаев.
                // Здесь мы просто сохраняем текущее значение, аналогично режиму хранения.
                default: begin
                    p_dout <= p_dout;
                end
            endcase
        end
    end

endmodule // Конец описания модуля universal_shift_reg
