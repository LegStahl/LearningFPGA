`timescale 1ns/1ns;
// Testbench - ??? ?????? ??? ?????? ?????-??????.
module adder_4bit_tb;
// 1. ????????? ?????????? ???? 'reg' ??? ?????? ????????
// ?? ????? ?????? ???????????? ?????????? (DUT).
reg [3:0] tb_a;
reg [3:0] tb_b;
reg tb_cin;
// 2. ????????? "???????" ???? 'wire' ??? ?????????? ????????
// ? ??????? ?????? DUT.
wire [3:0] tb_sum;
wire tb_cout;
// 3. ??????? ????????? (????????????) ???????????? ??????.
// ?????????, ??? ??? ?????? ???????? ?????? adder_4bit!
adder_4bit dut (
.a (tb_a),
.b (tb_b),
.cin (tb_cin),
.sum (tb_sum),
.cout (tb_cout)
);
// 4. ???? initial ????????? ???????? ????????????.
initial begin
// ? ????? ?????? ????????? ??????? ????????? ? ???????.
$display("?????\t A\t B\tCin | Cout\tSum");
$display("-------------------------------------------");
// ???? 1: 2 + 5 + 0 = 7
tb_a = 4'd2; tb_b = 4'd5; tb_cin = 1'b0;
#100; // ???? 10 ??????????, ????? ??????? ?????????.
// ???? 2: 9 + 1 + 0 = 10
tb_a = 4'd9; tb_b = 4'd1; tb_cin = 1'b0;
#100; // ???? ??? 10 ??.
// ???? 3: 15 + 1 + 0 = 16 (???????? ????????)
tb_a = 4'd15; tb_b = 4'd1; tb_cin = 1'b0;
#100;
// ???? 4: 8 + 8 + 1 = 17 (???????? ? ??????? ?????????)
tb_a = 4'd8; tb_b = 4'd8; tb_cin = 1'b1;
#100;
// ????????? ????????? ????? 10 ??.
#100 $finish;
end
// 5. (???????????) ???? $monitor ??? ???????? ??????.
initial begin
$monitor("%0t ns\t %d\t %d\t %b | %b\t\t%d", $time, tb_a, tb_b, tb_cin, tb_cout,
tb_sum);
end
endmodule
